//-------------------------------------------------------------------------------------------------
module ram
//-------------------------------------------------------------------------------------------------
#
(
	parameter KB = 0,
	parameter DW = 8
)
(
	input  wire                      clock,
	input  wire                      ce,
	input  wire                      we,
	input  wire[             DW-1:0] d,
	output reg [             DW-1:0] q,
	input  wire[$clog2(KB*1024)-1:0] a
);
//-------------------------------------------------------------------------------------------------

reg[DW-1:0] ram[(KB*1024)-1:0];

always @(posedge clock) if(ce) if(!we) ram[a] <= d; else q <= ram[a];

//-------------------------------------------------------------------------------------------------
endmodule
//-------------------------------------------------------------------------------------------------
