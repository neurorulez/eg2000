-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bab",
     9 => x"bc080b0b",
    10 => x"0babc008",
    11 => x"0b0b0bab",
    12 => x"c4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"abc40c0b",
    16 => x"0b0babc0",
    17 => x"0c0b0b0b",
    18 => x"abbc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0ba78c",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"abbc70b0",
    57 => x"e0278b38",
    58 => x"80717084",
    59 => x"05530c81",
    60 => x"e2048c51",
    61 => x"88e20402",
    62 => x"fc050df8",
    63 => x"80518f0b",
    64 => x"abcc0c9f",
    65 => x"0babd00c",
    66 => x"a0717081",
    67 => x"055334ab",
    68 => x"d008ff05",
    69 => x"abd00cab",
    70 => x"d0088025",
    71 => x"eb38abcc",
    72 => x"08ff05ab",
    73 => x"cc0cabcc",
    74 => x"088025d7",
    75 => x"38800bab",
    76 => x"d00c800b",
    77 => x"abcc0c02",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"abcc0825",
    97 => x"8f3882bc",
    98 => x"2dabcc08",
    99 => x"ff05abcc",
   100 => x"0c82fe04",
   101 => x"abcc08ab",
   102 => x"d0085351",
   103 => x"728a2e09",
   104 => x"8106b738",
   105 => x"7151719f",
   106 => x"24a038ab",
   107 => x"cc08a029",
   108 => x"11f88011",
   109 => x"5151a071",
   110 => x"34abd008",
   111 => x"8105abd0",
   112 => x"0cabd008",
   113 => x"519f7125",
   114 => x"e238800b",
   115 => x"abd00cab",
   116 => x"cc088105",
   117 => x"abcc0c83",
   118 => x"ee0470a0",
   119 => x"2912f880",
   120 => x"11515172",
   121 => x"7134abd0",
   122 => x"088105ab",
   123 => x"d00cabd0",
   124 => x"08a02e09",
   125 => x"81068e38",
   126 => x"800babd0",
   127 => x"0cabcc08",
   128 => x"8105abcc",
   129 => x"0c028c05",
   130 => x"0d0402e8",
   131 => x"050d7779",
   132 => x"5656880b",
   133 => x"fc167771",
   134 => x"2c8f0654",
   135 => x"52548053",
   136 => x"72722595",
   137 => x"387153fb",
   138 => x"e0145187",
   139 => x"71348114",
   140 => x"ff145454",
   141 => x"72f13871",
   142 => x"53f91576",
   143 => x"712c8706",
   144 => x"53517180",
   145 => x"2e8b38fb",
   146 => x"e0145171",
   147 => x"71348114",
   148 => x"54728e24",
   149 => x"95388f73",
   150 => x"3153fbe0",
   151 => x"1451a071",
   152 => x"348114ff",
   153 => x"14545472",
   154 => x"f1380298",
   155 => x"050d0402",
   156 => x"ec050d80",
   157 => x"0babd40c",
   158 => x"f68c08f6",
   159 => x"90087188",
   160 => x"2c565481",
   161 => x"ff065273",
   162 => x"72258838",
   163 => x"7154820b",
   164 => x"abd40c72",
   165 => x"882c7381",
   166 => x"ff065455",
   167 => x"7473258b",
   168 => x"3872abd4",
   169 => x"088407ab",
   170 => x"d40c5573",
   171 => x"842b86a0",
   172 => x"71258371",
   173 => x"31700b0b",
   174 => x"0ba9ec0c",
   175 => x"81712bff",
   176 => x"05f6880c",
   177 => x"fdfc13ff",
   178 => x"122c7888",
   179 => x"29ff9405",
   180 => x"70812cab",
   181 => x"d4085258",
   182 => x"52555152",
   183 => x"5476802e",
   184 => x"85387081",
   185 => x"075170f6",
   186 => x"940c7109",
   187 => x"8105f680",
   188 => x"0c720981",
   189 => x"05f6840c",
   190 => x"0294050d",
   191 => x"0402f405",
   192 => x"0d745372",
   193 => x"70810554",
   194 => x"80f52d52",
   195 => x"71802e89",
   196 => x"38715182",
   197 => x"f82d8683",
   198 => x"04810bab",
   199 => x"bc0c028c",
   200 => x"050d0402",
   201 => x"fc050d81",
   202 => x"808051c0",
   203 => x"115170fb",
   204 => x"38028405",
   205 => x"0d0402fc",
   206 => x"050d84bf",
   207 => x"5186a32d",
   208 => x"ff115170",
   209 => x"8025f638",
   210 => x"0284050d",
   211 => x"0402fc05",
   212 => x"0dec5183",
   213 => x"710c86a3",
   214 => x"2d82710c",
   215 => x"0284050d",
   216 => x"0402fc05",
   217 => x"0dec5192",
   218 => x"710c86a3",
   219 => x"2d82710c",
   220 => x"0284050d",
   221 => x"0402d005",
   222 => x"0d7d5480",
   223 => x"5ba40bec",
   224 => x"0c7352ab",
   225 => x"d851a3df",
   226 => x"2dabbc08",
   227 => x"7b2e81ab",
   228 => x"38abdc08",
   229 => x"70f80c89",
   230 => x"1580f52d",
   231 => x"8a1680f5",
   232 => x"2d718280",
   233 => x"29058817",
   234 => x"80f52d70",
   235 => x"84808029",
   236 => x"12f40c7e",
   237 => x"ff155c5e",
   238 => x"57555658",
   239 => x"767b2e8b",
   240 => x"38811a77",
   241 => x"812a585a",
   242 => x"76f738f7",
   243 => x"1a5a815b",
   244 => x"80782580",
   245 => x"e6387952",
   246 => x"7651848a",
   247 => x"2daca452",
   248 => x"abd851a6",
   249 => x"952dabbc",
   250 => x"08802eb8",
   251 => x"38aca45c",
   252 => x"83fc597b",
   253 => x"7084055d",
   254 => x"087081ff",
   255 => x"0671882a",
   256 => x"7081ff06",
   257 => x"73902a70",
   258 => x"81ff0675",
   259 => x"982ae80c",
   260 => x"e80c58e8",
   261 => x"0c57e80c",
   262 => x"fc1a5a53",
   263 => x"788025d3",
   264 => x"3888ab04",
   265 => x"abbc085b",
   266 => x"848058ab",
   267 => x"d851a5e8",
   268 => x"2dfc8018",
   269 => x"81185858",
   270 => x"87d00486",
   271 => x"b62d840b",
   272 => x"ec0c7a80",
   273 => x"2e8d38a9",
   274 => x"f0518eef",
   275 => x"2d8cf22d",
   276 => x"88d904aa",
   277 => x"c8518eef",
   278 => x"2d7aabbc",
   279 => x"0c02b005",
   280 => x"0d0402f4",
   281 => x"050d840b",
   282 => x"ec0c8cda",
   283 => x"2d89c42d",
   284 => x"81f72d9d",
   285 => x"ae2dabbc",
   286 => x"08802eb3",
   287 => x"3886f551",
   288 => x"a7872da9",
   289 => x"f0518eef",
   290 => x"2d8cf22d",
   291 => x"89d02d8e",
   292 => x"ff2daa9c",
   293 => x"0b80f52d",
   294 => x"70822b8c",
   295 => x"06fc0c53",
   296 => x"8652abbc",
   297 => x"08833884",
   298 => x"5271ec0c",
   299 => x"898c0480",
   300 => x"0babbc0c",
   301 => x"028c050d",
   302 => x"0471980c",
   303 => x"04ffb008",
   304 => x"abbc0c04",
   305 => x"810bffb0",
   306 => x"0c04800b",
   307 => x"ffb00c04",
   308 => x"02f4050d",
   309 => x"8ad204ab",
   310 => x"bc0881f0",
   311 => x"2e098106",
   312 => x"8938810b",
   313 => x"abac0c8a",
   314 => x"d204abbc",
   315 => x"0881e02e",
   316 => x"09810689",
   317 => x"38810bab",
   318 => x"b00c8ad2",
   319 => x"04abbc08",
   320 => x"52abb008",
   321 => x"802e8838",
   322 => x"abbc0881",
   323 => x"80055271",
   324 => x"842c728f",
   325 => x"065353ab",
   326 => x"ac08802e",
   327 => x"99387284",
   328 => x"29aaec05",
   329 => x"72138171",
   330 => x"2b700973",
   331 => x"0806730c",
   332 => x"5153538a",
   333 => x"c8047284",
   334 => x"29aaec05",
   335 => x"72138371",
   336 => x"2b720807",
   337 => x"720c5353",
   338 => x"800babb0",
   339 => x"0c800bab",
   340 => x"ac0cabe4",
   341 => x"518bd32d",
   342 => x"abbc08ff",
   343 => x"24fef838",
   344 => x"800babbc",
   345 => x"0c028c05",
   346 => x"0d0402f8",
   347 => x"050daaec",
   348 => x"528f5180",
   349 => x"72708405",
   350 => x"540cff11",
   351 => x"51708025",
   352 => x"f2380288",
   353 => x"050d0402",
   354 => x"f0050d75",
   355 => x"5189ca2d",
   356 => x"70822cfc",
   357 => x"06aaec11",
   358 => x"72109e06",
   359 => x"71087072",
   360 => x"2a708306",
   361 => x"82742b70",
   362 => x"09740676",
   363 => x"0c545156",
   364 => x"57535153",
   365 => x"89c42d71",
   366 => x"abbc0c02",
   367 => x"90050d04",
   368 => x"02fc050d",
   369 => x"72518071",
   370 => x"0c800b84",
   371 => x"120c0284",
   372 => x"050d0402",
   373 => x"f0050d75",
   374 => x"70088412",
   375 => x"08535353",
   376 => x"ff547171",
   377 => x"2ea83889",
   378 => x"ca2d8413",
   379 => x"08708429",
   380 => x"14881170",
   381 => x"087081ff",
   382 => x"06841808",
   383 => x"81118706",
   384 => x"841a0c53",
   385 => x"51555151",
   386 => x"5189c42d",
   387 => x"715473ab",
   388 => x"bc0c0290",
   389 => x"050d0402",
   390 => x"f8050d89",
   391 => x"ca2de008",
   392 => x"708b2a70",
   393 => x"81065152",
   394 => x"5270802e",
   395 => x"9d38abe4",
   396 => x"08708429",
   397 => x"abec0573",
   398 => x"81ff0671",
   399 => x"0c5151ab",
   400 => x"e4088111",
   401 => x"8706abe4",
   402 => x"0c51800b",
   403 => x"ac8c0c89",
   404 => x"bd2d89c4",
   405 => x"2d028805",
   406 => x"0d0402fc",
   407 => x"050dabe4",
   408 => x"518bc02d",
   409 => x"8aea2d8c",
   410 => x"975189b9",
   411 => x"2d028405",
   412 => x"0d0402fc",
   413 => x"050d8cfc",
   414 => x"0489d02d",
   415 => x"80f6518b",
   416 => x"872dabbc",
   417 => x"08f33880",
   418 => x"da518b87",
   419 => x"2dabbc08",
   420 => x"e838abbc",
   421 => x"08abb80c",
   422 => x"abbc0851",
   423 => x"84ef2d02",
   424 => x"84050d04",
   425 => x"02ec050d",
   426 => x"76548052",
   427 => x"870b8815",
   428 => x"80f52d56",
   429 => x"53747224",
   430 => x"8338a053",
   431 => x"725182f8",
   432 => x"2d81128b",
   433 => x"1580f52d",
   434 => x"54527272",
   435 => x"25de3802",
   436 => x"94050d04",
   437 => x"02f0050d",
   438 => x"ac900854",
   439 => x"81f72d80",
   440 => x"0bac940c",
   441 => x"7308802e",
   442 => x"81803882",
   443 => x"0babd00c",
   444 => x"ac94088f",
   445 => x"06abcc0c",
   446 => x"73085271",
   447 => x"832e9638",
   448 => x"71832689",
   449 => x"3871812e",
   450 => x"af388ed5",
   451 => x"0471852e",
   452 => x"9f388ed5",
   453 => x"04881480",
   454 => x"f52d8415",
   455 => x"08a8c053",
   456 => x"545285fd",
   457 => x"2d718429",
   458 => x"13700852",
   459 => x"528ed904",
   460 => x"73518da4",
   461 => x"2d8ed504",
   462 => x"abb40888",
   463 => x"15082c70",
   464 => x"81065152",
   465 => x"71802e87",
   466 => x"38a8c451",
   467 => x"8ed204a8",
   468 => x"c85185fd",
   469 => x"2d841408",
   470 => x"5185fd2d",
   471 => x"ac940881",
   472 => x"05ac940c",
   473 => x"8c14548d",
   474 => x"e4040290",
   475 => x"050d0471",
   476 => x"ac900c8d",
   477 => x"d42dac94",
   478 => x"08ff05ac",
   479 => x"980c0402",
   480 => x"e8050dac",
   481 => x"9008ac9c",
   482 => x"08575587",
   483 => x"518b872d",
   484 => x"abbc0881",
   485 => x"2a708106",
   486 => x"51527180",
   487 => x"2ea0388f",
   488 => x"a50489d0",
   489 => x"2d87518b",
   490 => x"872dabbc",
   491 => x"08f438ab",
   492 => x"b8088132",
   493 => x"70abb80c",
   494 => x"70525284",
   495 => x"ef2d80fe",
   496 => x"518b872d",
   497 => x"abbc0880",
   498 => x"2ea638ab",
   499 => x"b808802e",
   500 => x"9138800b",
   501 => x"abb80c80",
   502 => x"5184ef2d",
   503 => x"8fe20489",
   504 => x"d02d80fe",
   505 => x"518b872d",
   506 => x"abbc08f3",
   507 => x"3886e12d",
   508 => x"abb80890",
   509 => x"3881fd51",
   510 => x"8b872d81",
   511 => x"fa518b87",
   512 => x"2d95b504",
   513 => x"81f5518b",
   514 => x"872dabbc",
   515 => x"08812a70",
   516 => x"81065152",
   517 => x"71802eaf",
   518 => x"38ac9808",
   519 => x"5271802e",
   520 => x"8938ff12",
   521 => x"ac980c90",
   522 => x"c704ac94",
   523 => x"0810ac94",
   524 => x"08057084",
   525 => x"29165152",
   526 => x"88120880",
   527 => x"2e8938ff",
   528 => x"51881208",
   529 => x"52712d81",
   530 => x"f2518b87",
   531 => x"2dabbc08",
   532 => x"812a7081",
   533 => x"06515271",
   534 => x"802eb138",
   535 => x"ac9408ff",
   536 => x"11ac9808",
   537 => x"56535373",
   538 => x"72258938",
   539 => x"8114ac98",
   540 => x"0c918c04",
   541 => x"72101370",
   542 => x"84291651",
   543 => x"52881208",
   544 => x"802e8938",
   545 => x"fe518812",
   546 => x"0852712d",
   547 => x"81fd518b",
   548 => x"872dabbc",
   549 => x"08812a70",
   550 => x"81065152",
   551 => x"71802ead",
   552 => x"38ac9808",
   553 => x"802e8938",
   554 => x"800bac98",
   555 => x"0c91cd04",
   556 => x"ac940810",
   557 => x"ac940805",
   558 => x"70842916",
   559 => x"51528812",
   560 => x"08802e89",
   561 => x"38fd5188",
   562 => x"12085271",
   563 => x"2d81fa51",
   564 => x"8b872dab",
   565 => x"bc08812a",
   566 => x"70810651",
   567 => x"5271802e",
   568 => x"ae38ac94",
   569 => x"08ff1154",
   570 => x"52ac9808",
   571 => x"73258838",
   572 => x"72ac980c",
   573 => x"928f0471",
   574 => x"10127084",
   575 => x"29165152",
   576 => x"88120880",
   577 => x"2e8938fc",
   578 => x"51881208",
   579 => x"52712dac",
   580 => x"98087053",
   581 => x"5473802e",
   582 => x"8a388c15",
   583 => x"ff155555",
   584 => x"92950482",
   585 => x"0babd00c",
   586 => x"718f06ab",
   587 => x"cc0c81eb",
   588 => x"518b872d",
   589 => x"abbc0881",
   590 => x"2a708106",
   591 => x"51527180",
   592 => x"2ead3874",
   593 => x"08852e09",
   594 => x"8106a438",
   595 => x"881580f5",
   596 => x"2dff0552",
   597 => x"71881681",
   598 => x"b72d7198",
   599 => x"2b527180",
   600 => x"25883880",
   601 => x"0b881681",
   602 => x"b72d7451",
   603 => x"8da42d81",
   604 => x"f4518b87",
   605 => x"2dabbc08",
   606 => x"812a7081",
   607 => x"06515271",
   608 => x"802eb338",
   609 => x"7408852e",
   610 => x"098106aa",
   611 => x"38881580",
   612 => x"f52d8105",
   613 => x"52718816",
   614 => x"81b72d71",
   615 => x"81ff068b",
   616 => x"1680f52d",
   617 => x"54527272",
   618 => x"27873872",
   619 => x"881681b7",
   620 => x"2d74518d",
   621 => x"a42d80da",
   622 => x"518b872d",
   623 => x"abbc0881",
   624 => x"2a708106",
   625 => x"51527180",
   626 => x"2e81a638",
   627 => x"ac9008ac",
   628 => x"98085553",
   629 => x"73802e8a",
   630 => x"388c13ff",
   631 => x"15555393",
   632 => x"d4047208",
   633 => x"5271822e",
   634 => x"a6387182",
   635 => x"26893871",
   636 => x"812ea938",
   637 => x"94f10471",
   638 => x"832eb138",
   639 => x"71842e09",
   640 => x"810680ed",
   641 => x"38881308",
   642 => x"518eef2d",
   643 => x"94f104ac",
   644 => x"98085188",
   645 => x"13085271",
   646 => x"2d94f104",
   647 => x"810b8814",
   648 => x"082babb4",
   649 => x"0832abb4",
   650 => x"0c94c704",
   651 => x"881380f5",
   652 => x"2d81058b",
   653 => x"1480f52d",
   654 => x"53547174",
   655 => x"24833880",
   656 => x"54738814",
   657 => x"81b72d8d",
   658 => x"d42d94f1",
   659 => x"04750880",
   660 => x"2ea23875",
   661 => x"08518b87",
   662 => x"2dabbc08",
   663 => x"81065271",
   664 => x"802e8b38",
   665 => x"ac980851",
   666 => x"84160852",
   667 => x"712d8816",
   668 => x"5675da38",
   669 => x"8054800b",
   670 => x"abd00c73",
   671 => x"8f06abcc",
   672 => x"0ca05273",
   673 => x"ac98082e",
   674 => x"09810698",
   675 => x"38ac9408",
   676 => x"ff057432",
   677 => x"70098105",
   678 => x"7072079f",
   679 => x"2a917131",
   680 => x"51515353",
   681 => x"715182f8",
   682 => x"2d811454",
   683 => x"8e7425c6",
   684 => x"38abb808",
   685 => x"5271abbc",
   686 => x"0c029805",
   687 => x"0d0402f4",
   688 => x"050dd452",
   689 => x"81ff720c",
   690 => x"71085381",
   691 => x"ff720c72",
   692 => x"882b83fe",
   693 => x"80067208",
   694 => x"7081ff06",
   695 => x"51525381",
   696 => x"ff720c72",
   697 => x"7107882b",
   698 => x"72087081",
   699 => x"ff065152",
   700 => x"5381ff72",
   701 => x"0c727107",
   702 => x"882b7208",
   703 => x"7081ff06",
   704 => x"7207abbc",
   705 => x"0c525302",
   706 => x"8c050d04",
   707 => x"02f4050d",
   708 => x"74767181",
   709 => x"ff06d40c",
   710 => x"5353aca0",
   711 => x"08853871",
   712 => x"892b5271",
   713 => x"982ad40c",
   714 => x"71902a70",
   715 => x"81ff06d4",
   716 => x"0c517188",
   717 => x"2a7081ff",
   718 => x"06d40c51",
   719 => x"7181ff06",
   720 => x"d40c7290",
   721 => x"2a7081ff",
   722 => x"06d40c51",
   723 => x"d4087081",
   724 => x"ff065151",
   725 => x"82b8bf52",
   726 => x"7081ff2e",
   727 => x"09810694",
   728 => x"3881ff0b",
   729 => x"d40cd408",
   730 => x"7081ff06",
   731 => x"ff145451",
   732 => x"5171e538",
   733 => x"70abbc0c",
   734 => x"028c050d",
   735 => x"0402fc05",
   736 => x"0d81c751",
   737 => x"81ff0bd4",
   738 => x"0cff1151",
   739 => x"708025f4",
   740 => x"38028405",
   741 => x"0d0402f4",
   742 => x"050d81ff",
   743 => x"0bd40c93",
   744 => x"53805287",
   745 => x"fc80c151",
   746 => x"968c2dab",
   747 => x"bc088b38",
   748 => x"81ff0bd4",
   749 => x"0c815397",
   750 => x"c30496fd",
   751 => x"2dff1353",
   752 => x"72df3872",
   753 => x"abbc0c02",
   754 => x"8c050d04",
   755 => x"02ec050d",
   756 => x"810baca0",
   757 => x"0c8454d0",
   758 => x"08708f2a",
   759 => x"70810651",
   760 => x"515372f3",
   761 => x"3872d00c",
   762 => x"96fd2da8",
   763 => x"cc5185fd",
   764 => x"2dd00870",
   765 => x"8f2a7081",
   766 => x"06515153",
   767 => x"72f33881",
   768 => x"0bd00cb1",
   769 => x"53805284",
   770 => x"d480c051",
   771 => x"968c2dab",
   772 => x"bc08812e",
   773 => x"93387282",
   774 => x"2ebd38ff",
   775 => x"135372e5",
   776 => x"38ff1454",
   777 => x"73ffb038",
   778 => x"96fd2d83",
   779 => x"aa52849c",
   780 => x"80c85196",
   781 => x"8c2dabbc",
   782 => x"08812e09",
   783 => x"81069238",
   784 => x"95be2dab",
   785 => x"bc0883ff",
   786 => x"ff065372",
   787 => x"83aa2e9d",
   788 => x"3897962d",
   789 => x"98e804a8",
   790 => x"d85185fd",
   791 => x"2d80539a",
   792 => x"b604a8f0",
   793 => x"5185fd2d",
   794 => x"80549a88",
   795 => x"0481ff0b",
   796 => x"d40cb154",
   797 => x"96fd2d8f",
   798 => x"cf538052",
   799 => x"87fc80f7",
   800 => x"51968c2d",
   801 => x"abbc0855",
   802 => x"abbc0881",
   803 => x"2e098106",
   804 => x"9b3881ff",
   805 => x"0bd40c82",
   806 => x"0a52849c",
   807 => x"80e95196",
   808 => x"8c2dabbc",
   809 => x"08802e8d",
   810 => x"3896fd2d",
   811 => x"ff135372",
   812 => x"c93899fb",
   813 => x"0481ff0b",
   814 => x"d40cabbc",
   815 => x"085287fc",
   816 => x"80fa5196",
   817 => x"8c2dabbc",
   818 => x"08b13881",
   819 => x"ff0bd40c",
   820 => x"d4085381",
   821 => x"ff0bd40c",
   822 => x"81ff0bd4",
   823 => x"0c81ff0b",
   824 => x"d40c81ff",
   825 => x"0bd40c72",
   826 => x"862a7081",
   827 => x"06765651",
   828 => x"53729538",
   829 => x"abbc0854",
   830 => x"9a880473",
   831 => x"822efee2",
   832 => x"38ff1454",
   833 => x"73feed38",
   834 => x"73aca00c",
   835 => x"738b3881",
   836 => x"5287fc80",
   837 => x"d051968c",
   838 => x"2d81ff0b",
   839 => x"d40cd008",
   840 => x"708f2a70",
   841 => x"81065151",
   842 => x"5372f338",
   843 => x"72d00c81",
   844 => x"ff0bd40c",
   845 => x"815372ab",
   846 => x"bc0c0294",
   847 => x"050d0402",
   848 => x"e8050d78",
   849 => x"55805681",
   850 => x"ff0bd40c",
   851 => x"d008708f",
   852 => x"2a708106",
   853 => x"51515372",
   854 => x"f3388281",
   855 => x"0bd00c81",
   856 => x"ff0bd40c",
   857 => x"775287fc",
   858 => x"80d15196",
   859 => x"8c2d80db",
   860 => x"c6df54ab",
   861 => x"bc08802e",
   862 => x"8a38a990",
   863 => x"5185fd2d",
   864 => x"9bd60481",
   865 => x"ff0bd40c",
   866 => x"d4087081",
   867 => x"ff065153",
   868 => x"7281fe2e",
   869 => x"0981069d",
   870 => x"3880ff53",
   871 => x"95be2dab",
   872 => x"bc087570",
   873 => x"8405570c",
   874 => x"ff135372",
   875 => x"8025ed38",
   876 => x"81569bbb",
   877 => x"04ff1454",
   878 => x"73c93881",
   879 => x"ff0bd40c",
   880 => x"81ff0bd4",
   881 => x"0cd00870",
   882 => x"8f2a7081",
   883 => x"06515153",
   884 => x"72f33872",
   885 => x"d00c75ab",
   886 => x"bc0c0298",
   887 => x"050d0402",
   888 => x"e8050d77",
   889 => x"797b5855",
   890 => x"55805372",
   891 => x"7625a338",
   892 => x"74708105",
   893 => x"5680f52d",
   894 => x"74708105",
   895 => x"5680f52d",
   896 => x"52527171",
   897 => x"2e863881",
   898 => x"519c9404",
   899 => x"8113539b",
   900 => x"eb048051",
   901 => x"70abbc0c",
   902 => x"0298050d",
   903 => x"0402ec05",
   904 => x"0d765574",
   905 => x"802ebb38",
   906 => x"9a1580e0",
   907 => x"2d51a6eb",
   908 => x"2dabbc08",
   909 => x"abbc08b0",
   910 => x"d00cabbc",
   911 => x"085454b0",
   912 => x"ac08802e",
   913 => x"99389415",
   914 => x"80e02d51",
   915 => x"a6eb2dab",
   916 => x"bc08902b",
   917 => x"83fff00a",
   918 => x"06707507",
   919 => x"515372b0",
   920 => x"d00cb0d0",
   921 => x"08537280",
   922 => x"2e9938b0",
   923 => x"a408fe14",
   924 => x"7129b0b8",
   925 => x"0805b0d4",
   926 => x"0c70842b",
   927 => x"b0b00c54",
   928 => x"9da904b0",
   929 => x"bc08b0d0",
   930 => x"0cb0c008",
   931 => x"b0d40cb0",
   932 => x"ac08802e",
   933 => x"8a38b0a4",
   934 => x"08842b53",
   935 => x"9da504b0",
   936 => x"c408842b",
   937 => x"5372b0b0",
   938 => x"0c029405",
   939 => x"0d0402d8",
   940 => x"050d800b",
   941 => x"b0ac0c84",
   942 => x"5497cc2d",
   943 => x"abbc0880",
   944 => x"2e9538ac",
   945 => x"a4528051",
   946 => x"9abf2dab",
   947 => x"bc08802e",
   948 => x"8638fe54",
   949 => x"9ddf04ff",
   950 => x"14547380",
   951 => x"24db3873",
   952 => x"8c38a9a0",
   953 => x"5185fd2d",
   954 => x"7355a2e8",
   955 => x"04805681",
   956 => x"0bb0d80c",
   957 => x"8853a9b4",
   958 => x"52acda51",
   959 => x"9bdf2dab",
   960 => x"bc08762e",
   961 => x"09810687",
   962 => x"38abbc08",
   963 => x"b0d80c88",
   964 => x"53a9c052",
   965 => x"acf6519b",
   966 => x"df2dabbc",
   967 => x"088738ab",
   968 => x"bc08b0d8",
   969 => x"0cb0d808",
   970 => x"802e80f6",
   971 => x"38afea0b",
   972 => x"80f52daf",
   973 => x"eb0b80f5",
   974 => x"2d71982b",
   975 => x"71902b07",
   976 => x"afec0b80",
   977 => x"f52d7088",
   978 => x"2b7207af",
   979 => x"ed0b80f5",
   980 => x"2d7107b0",
   981 => x"a20b80f5",
   982 => x"2db0a30b",
   983 => x"80f52d71",
   984 => x"882b0753",
   985 => x"5f54525a",
   986 => x"56575573",
   987 => x"81abaa2e",
   988 => x"0981068d",
   989 => x"387551a6",
   990 => x"bb2dabbc",
   991 => x"08569f8e",
   992 => x"047382d4",
   993 => x"d52e8738",
   994 => x"a9cc519f",
   995 => x"cf04aca4",
   996 => x"5275519a",
   997 => x"bf2dabbc",
   998 => x"0855abbc",
   999 => x"08802e83",
  1000 => x"c7388853",
  1001 => x"a9c052ac",
  1002 => x"f6519bdf",
  1003 => x"2dabbc08",
  1004 => x"8938810b",
  1005 => x"b0ac0c9f",
  1006 => x"d5048853",
  1007 => x"a9b452ac",
  1008 => x"da519bdf",
  1009 => x"2dabbc08",
  1010 => x"802e8a38",
  1011 => x"a9e05185",
  1012 => x"fd2da0af",
  1013 => x"04b0a20b",
  1014 => x"80f52d54",
  1015 => x"7380d52e",
  1016 => x"09810680",
  1017 => x"ca38b0a3",
  1018 => x"0b80f52d",
  1019 => x"547381aa",
  1020 => x"2e098106",
  1021 => x"ba38800b",
  1022 => x"aca40b80",
  1023 => x"f52d5654",
  1024 => x"7481e92e",
  1025 => x"83388154",
  1026 => x"7481eb2e",
  1027 => x"8c388055",
  1028 => x"73752e09",
  1029 => x"810682d0",
  1030 => x"38acaf0b",
  1031 => x"80f52d55",
  1032 => x"748d38ac",
  1033 => x"b00b80f5",
  1034 => x"2d547382",
  1035 => x"2e863880",
  1036 => x"55a2e804",
  1037 => x"acb10b80",
  1038 => x"f52d70b0",
  1039 => x"a40cff05",
  1040 => x"b0a80cac",
  1041 => x"b20b80f5",
  1042 => x"2dacb30b",
  1043 => x"80f52d58",
  1044 => x"76057782",
  1045 => x"80290570",
  1046 => x"b0b40cac",
  1047 => x"b40b80f5",
  1048 => x"2d70b0c8",
  1049 => x"0cb0ac08",
  1050 => x"59575876",
  1051 => x"802e81a3",
  1052 => x"388853a9",
  1053 => x"c052acf6",
  1054 => x"519bdf2d",
  1055 => x"abbc0881",
  1056 => x"e738b0a4",
  1057 => x"0870842b",
  1058 => x"b0b00c70",
  1059 => x"b0c40cac",
  1060 => x"c90b80f5",
  1061 => x"2dacc80b",
  1062 => x"80f52d71",
  1063 => x"82802905",
  1064 => x"acca0b80",
  1065 => x"f52d7084",
  1066 => x"80802912",
  1067 => x"accb0b80",
  1068 => x"f52d7081",
  1069 => x"800a2912",
  1070 => x"70b0cc0c",
  1071 => x"b0c80871",
  1072 => x"29b0b408",
  1073 => x"0570b0b8",
  1074 => x"0cacd10b",
  1075 => x"80f52dac",
  1076 => x"d00b80f5",
  1077 => x"2d718280",
  1078 => x"2905acd2",
  1079 => x"0b80f52d",
  1080 => x"70848080",
  1081 => x"2912acd3",
  1082 => x"0b80f52d",
  1083 => x"70982b81",
  1084 => x"f00a0672",
  1085 => x"0570b0bc",
  1086 => x"0cfe117e",
  1087 => x"297705b0",
  1088 => x"c00c5259",
  1089 => x"5243545e",
  1090 => x"51525952",
  1091 => x"5d575957",
  1092 => x"a2e104ac",
  1093 => x"b60b80f5",
  1094 => x"2dacb50b",
  1095 => x"80f52d71",
  1096 => x"82802905",
  1097 => x"70b0b00c",
  1098 => x"70a02983",
  1099 => x"ff057089",
  1100 => x"2a70b0c4",
  1101 => x"0cacbb0b",
  1102 => x"80f52dac",
  1103 => x"ba0b80f5",
  1104 => x"2d718280",
  1105 => x"290570b0",
  1106 => x"cc0c7b71",
  1107 => x"291e70b0",
  1108 => x"c00c7db0",
  1109 => x"bc0c7305",
  1110 => x"b0b80c55",
  1111 => x"5e515155",
  1112 => x"5580519c",
  1113 => x"9d2d8155",
  1114 => x"74abbc0c",
  1115 => x"02a8050d",
  1116 => x"0402ec05",
  1117 => x"0d767087",
  1118 => x"2c7180ff",
  1119 => x"06555654",
  1120 => x"b0ac088a",
  1121 => x"3873882c",
  1122 => x"7481ff06",
  1123 => x"5455aca4",
  1124 => x"52b0b408",
  1125 => x"15519abf",
  1126 => x"2dabbc08",
  1127 => x"54abbc08",
  1128 => x"802eb338",
  1129 => x"b0ac0880",
  1130 => x"2e983872",
  1131 => x"8429aca4",
  1132 => x"05700852",
  1133 => x"53a6bb2d",
  1134 => x"abbc08f0",
  1135 => x"0a0653a3",
  1136 => x"d4047210",
  1137 => x"aca40570",
  1138 => x"80e02d52",
  1139 => x"53a6eb2d",
  1140 => x"abbc0853",
  1141 => x"725473ab",
  1142 => x"bc0c0294",
  1143 => x"050d0402",
  1144 => x"cc050d7e",
  1145 => x"605e5a80",
  1146 => x"0bb0d008",
  1147 => x"b0d40859",
  1148 => x"5c568058",
  1149 => x"b0b00878",
  1150 => x"2e81ae38",
  1151 => x"778f06a0",
  1152 => x"17575473",
  1153 => x"8f38aca4",
  1154 => x"52765181",
  1155 => x"17579abf",
  1156 => x"2daca456",
  1157 => x"807680f5",
  1158 => x"2d565474",
  1159 => x"742e8338",
  1160 => x"81547481",
  1161 => x"e52e80f6",
  1162 => x"38817075",
  1163 => x"06555c73",
  1164 => x"802e80ea",
  1165 => x"388b1680",
  1166 => x"f52d9806",
  1167 => x"597880de",
  1168 => x"388b537c",
  1169 => x"5275519b",
  1170 => x"df2dabbc",
  1171 => x"0880cf38",
  1172 => x"9c160851",
  1173 => x"a6bb2dab",
  1174 => x"bc08841b",
  1175 => x"0c9a1680",
  1176 => x"e02d51a6",
  1177 => x"eb2dabbc",
  1178 => x"08abbc08",
  1179 => x"881c0cab",
  1180 => x"bc085555",
  1181 => x"b0ac0880",
  1182 => x"2e983894",
  1183 => x"1680e02d",
  1184 => x"51a6eb2d",
  1185 => x"abbc0890",
  1186 => x"2b83fff0",
  1187 => x"0a067016",
  1188 => x"51547388",
  1189 => x"1b0c787a",
  1190 => x"0c7b54a5",
  1191 => x"df048118",
  1192 => x"58b0b008",
  1193 => x"7826fed4",
  1194 => x"38b0ac08",
  1195 => x"802eae38",
  1196 => x"7a51a2f1",
  1197 => x"2dabbc08",
  1198 => x"abbc0880",
  1199 => x"fffffff8",
  1200 => x"06555b73",
  1201 => x"80ffffff",
  1202 => x"f82e9238",
  1203 => x"abbc08fe",
  1204 => x"05b0a408",
  1205 => x"29b0b808",
  1206 => x"0557a3f2",
  1207 => x"04805473",
  1208 => x"abbc0c02",
  1209 => x"b4050d04",
  1210 => x"02f4050d",
  1211 => x"74700881",
  1212 => x"05710c70",
  1213 => x"08b0a808",
  1214 => x"06535371",
  1215 => x"8e388813",
  1216 => x"0851a2f1",
  1217 => x"2dabbc08",
  1218 => x"88140c81",
  1219 => x"0babbc0c",
  1220 => x"028c050d",
  1221 => x"0402f005",
  1222 => x"0d758811",
  1223 => x"08fe05b0",
  1224 => x"a40829b0",
  1225 => x"b8081172",
  1226 => x"08b0a808",
  1227 => x"06057955",
  1228 => x"5354549a",
  1229 => x"bf2d0290",
  1230 => x"050d0402",
  1231 => x"f4050d74",
  1232 => x"70882a83",
  1233 => x"fe800670",
  1234 => x"72982a07",
  1235 => x"72882b87",
  1236 => x"fc808006",
  1237 => x"73982b81",
  1238 => x"f00a0671",
  1239 => x"730707ab",
  1240 => x"bc0c5651",
  1241 => x"5351028c",
  1242 => x"050d0402",
  1243 => x"f8050d02",
  1244 => x"8e0580f5",
  1245 => x"2d74882b",
  1246 => x"077083ff",
  1247 => x"ff06abbc",
  1248 => x"0c510288",
  1249 => x"050d0471",
  1250 => x"b0dc0c04",
  1251 => x"00ffffff",
  1252 => x"ff00ffff",
  1253 => x"ffff00ff",
  1254 => x"ffffff00",
  1255 => x"20202020",
  1256 => x"203d4547",
  1257 => x"32303030",
  1258 => x"3d202020",
  1259 => x"20200000",
  1260 => x"20202020",
  1261 => x"4e657572",
  1262 => x"6f52756c",
  1263 => x"657a2020",
  1264 => x"20200000",
  1265 => x"52657365",
  1266 => x"74000000",
  1267 => x"45786974",
  1268 => x"00000000",
  1269 => x"5363616e",
  1270 => x"646f7562",
  1271 => x"6c657246",
  1272 => x"78204e6f",
  1273 => x"6e650000",
  1274 => x"5363616e",
  1275 => x"646f7562",
  1276 => x"6c657246",
  1277 => x"78204851",
  1278 => x"32780000",
  1279 => x"5363616e",
  1280 => x"646f7562",
  1281 => x"6c657246",
  1282 => x"78204352",
  1283 => x"54203235",
  1284 => x"25000000",
  1285 => x"5363616e",
  1286 => x"646f7562",
  1287 => x"6c657246",
  1288 => x"78204352",
  1289 => x"54203530",
  1290 => x"25000000",
  1291 => x"43617267",
  1292 => x"61204661",
  1293 => x"6c6c6964",
  1294 => x"61000000",
  1295 => x"4f4b0000",
  1296 => x"16200000",
  1297 => x"14200000",
  1298 => x"15200000",
  1299 => x"53442069",
  1300 => x"6e69742e",
  1301 => x"2e2e0a00",
  1302 => x"53442063",
  1303 => x"61726420",
  1304 => x"72657365",
  1305 => x"74206661",
  1306 => x"696c6564",
  1307 => x"210a0000",
  1308 => x"53444843",
  1309 => x"20657272",
  1310 => x"6f72210a",
  1311 => x"00000000",
  1312 => x"57726974",
  1313 => x"65206661",
  1314 => x"696c6564",
  1315 => x"0a000000",
  1316 => x"52656164",
  1317 => x"20666169",
  1318 => x"6c65640a",
  1319 => x"00000000",
  1320 => x"43617264",
  1321 => x"20696e69",
  1322 => x"74206661",
  1323 => x"696c6564",
  1324 => x"0a000000",
  1325 => x"46415431",
  1326 => x"36202020",
  1327 => x"00000000",
  1328 => x"46415433",
  1329 => x"32202020",
  1330 => x"00000000",
  1331 => x"4e6f2070",
  1332 => x"61727469",
  1333 => x"74696f6e",
  1334 => x"20736967",
  1335 => x"0a000000",
  1336 => x"42616420",
  1337 => x"70617274",
  1338 => x"0a000000",
  1339 => x"00000002",
  1340 => x"00000002",
  1341 => x"0000139c",
  1342 => x"00000000",
  1343 => x"00000002",
  1344 => x"000013b0",
  1345 => x"00000000",
  1346 => x"00000002",
  1347 => x"000013c4",
  1348 => x"0000034d",
  1349 => x"00000003",
  1350 => x"00001538",
  1351 => x"00000004",
  1352 => x"00000002",
  1353 => x"000013cc",
  1354 => x"00000672",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"000013d4",
  1359 => x"000013e8",
  1360 => x"000013fc",
  1361 => x"00001414",
  1362 => x"00000004",
  1363 => x"0000142c",
  1364 => x"00001548",
  1365 => x"00000004",
  1366 => x"0000143c",
  1367 => x"000014f0",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

